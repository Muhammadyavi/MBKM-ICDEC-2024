magic
tech sky130A
magscale 1 2
timestamp 1729314602
<< nwell >>
rect 2785 535 4582 1641
<< pmos >>
rect 3027 1221 3057 1421
rect 3227 1221 3327 1421
rect 3499 1221 3599 1421
rect 3771 1221 3871 1421
rect 4043 1221 4143 1421
rect 4313 1221 4343 1421
rect 3027 785 3057 985
rect 3227 785 3327 985
rect 3499 785 3599 985
rect 3771 785 3871 985
rect 4043 785 4143 985
rect 4313 785 4343 985
<< pdiff >>
rect 2969 1409 3027 1421
rect 2969 1233 2981 1409
rect 3015 1233 3027 1409
rect 2969 1221 3027 1233
rect 3057 1409 3115 1421
rect 3057 1233 3069 1409
rect 3103 1233 3115 1409
rect 3057 1221 3115 1233
rect 3169 1409 3227 1421
rect 3169 1233 3181 1409
rect 3215 1233 3227 1409
rect 3169 1221 3227 1233
rect 3327 1409 3385 1421
rect 3327 1233 3339 1409
rect 3373 1233 3385 1409
rect 3327 1221 3385 1233
rect 3441 1409 3499 1421
rect 3441 1233 3453 1409
rect 3487 1233 3499 1409
rect 3441 1221 3499 1233
rect 3599 1409 3657 1421
rect 3599 1233 3611 1409
rect 3645 1233 3657 1409
rect 3599 1221 3657 1233
rect 3713 1409 3771 1421
rect 3713 1233 3725 1409
rect 3759 1233 3771 1409
rect 3713 1221 3771 1233
rect 3871 1409 3929 1421
rect 3871 1233 3883 1409
rect 3917 1233 3929 1409
rect 3871 1221 3929 1233
rect 3985 1409 4043 1421
rect 3985 1233 3997 1409
rect 4031 1233 4043 1409
rect 3985 1221 4043 1233
rect 4143 1409 4201 1421
rect 4143 1233 4155 1409
rect 4189 1233 4201 1409
rect 4143 1221 4201 1233
rect 4255 1409 4313 1421
rect 4255 1233 4267 1409
rect 4301 1233 4313 1409
rect 4255 1221 4313 1233
rect 4343 1409 4401 1421
rect 4343 1233 4355 1409
rect 4389 1233 4401 1409
rect 4343 1221 4401 1233
rect 2969 973 3027 985
rect 2969 797 2981 973
rect 3015 797 3027 973
rect 2969 785 3027 797
rect 3057 973 3115 985
rect 3057 797 3069 973
rect 3103 797 3115 973
rect 3057 785 3115 797
rect 3169 973 3227 985
rect 3169 797 3181 973
rect 3215 797 3227 973
rect 3169 785 3227 797
rect 3327 973 3385 985
rect 3327 797 3339 973
rect 3373 797 3385 973
rect 3327 785 3385 797
rect 3441 973 3499 985
rect 3441 797 3453 973
rect 3487 797 3499 973
rect 3441 785 3499 797
rect 3599 973 3657 985
rect 3599 797 3611 973
rect 3645 797 3657 973
rect 3599 785 3657 797
rect 3713 973 3771 985
rect 3713 797 3725 973
rect 3759 797 3771 973
rect 3713 785 3771 797
rect 3871 973 3929 985
rect 3871 797 3883 973
rect 3917 797 3929 973
rect 3871 785 3929 797
rect 3985 973 4043 985
rect 3985 797 3997 973
rect 4031 797 4043 973
rect 3985 785 4043 797
rect 4143 973 4201 985
rect 4143 797 4155 973
rect 4189 797 4201 973
rect 4143 785 4201 797
rect 4255 973 4313 985
rect 4255 797 4267 973
rect 4301 797 4313 973
rect 4255 785 4313 797
rect 4343 973 4401 985
rect 4343 797 4355 973
rect 4389 797 4401 973
rect 4343 785 4401 797
<< pdiffc >>
rect 2981 1233 3015 1409
rect 3069 1233 3103 1409
rect 3181 1233 3215 1409
rect 3339 1233 3373 1409
rect 3453 1233 3487 1409
rect 3611 1233 3645 1409
rect 3725 1233 3759 1409
rect 3883 1233 3917 1409
rect 3997 1233 4031 1409
rect 4155 1233 4189 1409
rect 4267 1233 4301 1409
rect 4355 1233 4389 1409
rect 2981 797 3015 973
rect 3069 797 3103 973
rect 3181 797 3215 973
rect 3339 797 3373 973
rect 3453 797 3487 973
rect 3611 797 3645 973
rect 3725 797 3759 973
rect 3883 797 3917 973
rect 3997 797 4031 973
rect 4155 797 4189 973
rect 4267 797 4301 973
rect 4355 797 4389 973
<< nsubdiff >>
rect 2821 1571 2881 1605
rect 4486 1571 4546 1605
rect 2821 1545 2855 1571
rect 4512 1545 4546 1571
rect 2821 605 2855 631
rect 4512 605 4546 631
rect 2821 571 2881 605
rect 4486 571 4546 605
<< nsubdiffcont >>
rect 2881 1571 4486 1605
rect 2821 631 2855 1545
rect 4512 631 4546 1545
rect 2881 571 4486 605
<< poly >>
rect 2965 1504 3057 1519
rect 2965 1470 2981 1504
rect 3015 1470 3057 1504
rect 2965 1451 3057 1470
rect 3027 1421 3057 1451
rect 3227 1508 3327 1518
rect 3499 1508 3599 1518
rect 3227 1502 3599 1508
rect 3227 1468 3243 1502
rect 3311 1468 3515 1502
rect 3583 1468 3599 1502
rect 3227 1462 3599 1468
rect 3227 1421 3327 1462
rect 3499 1421 3599 1462
rect 3771 1507 3871 1518
rect 4043 1507 4143 1518
rect 3771 1502 4143 1507
rect 3771 1468 3787 1502
rect 3855 1468 4059 1502
rect 4127 1468 4143 1502
rect 3771 1461 4143 1468
rect 3771 1421 3871 1461
rect 4043 1421 4143 1461
rect 4313 1503 4405 1518
rect 4313 1469 4355 1503
rect 4389 1469 4405 1503
rect 4313 1450 4405 1469
rect 4313 1421 4343 1450
rect 3027 1195 3057 1221
rect 3227 1181 3327 1221
rect 3499 1174 3599 1221
rect 3499 1140 3515 1174
rect 3583 1140 3599 1174
rect 3499 1124 3599 1140
rect 3771 1174 3871 1221
rect 4043 1183 4143 1221
rect 4313 1195 4343 1221
rect 3771 1140 3787 1174
rect 3855 1140 3871 1174
rect 3771 1124 3871 1140
rect 3499 1066 3599 1082
rect 3499 1032 3515 1066
rect 3583 1032 3599 1066
rect 3027 985 3057 1011
rect 3227 985 3327 1024
rect 3499 985 3599 1032
rect 3771 1066 3871 1082
rect 3771 1032 3787 1066
rect 3855 1032 3871 1066
rect 3771 985 3871 1032
rect 4043 985 4143 1026
rect 4313 985 4343 1011
rect 3027 745 3057 785
rect 2965 726 3057 745
rect 2965 692 2981 726
rect 3015 692 3057 726
rect 2965 677 3057 692
rect 3227 744 3327 785
rect 3499 744 3599 785
rect 3227 738 3599 744
rect 3227 704 3243 738
rect 3311 704 3515 738
rect 3583 704 3599 738
rect 3227 698 3599 704
rect 3227 688 3327 698
rect 3499 688 3599 698
rect 3771 744 3871 785
rect 4043 744 4143 785
rect 3771 738 4143 744
rect 3771 704 3787 738
rect 3855 704 4059 738
rect 4127 704 4143 738
rect 3771 698 4143 704
rect 3771 688 3871 698
rect 4043 688 4143 698
rect 4313 753 4343 785
rect 4313 734 4405 753
rect 4313 700 4355 734
rect 4389 700 4405 734
rect 4313 685 4405 700
<< polycont >>
rect 2981 1470 3015 1504
rect 3243 1468 3311 1502
rect 3515 1468 3583 1502
rect 3787 1468 3855 1502
rect 4059 1468 4127 1502
rect 4355 1469 4389 1503
rect 3515 1140 3583 1174
rect 3787 1140 3855 1174
rect 3515 1032 3583 1066
rect 3787 1032 3855 1066
rect 2981 692 3015 726
rect 3243 704 3311 738
rect 3515 704 3583 738
rect 3787 704 3855 738
rect 4059 704 4127 738
rect 4355 700 4389 734
<< locali >>
rect 2855 1571 2881 1605
rect 4486 1572 4512 1605
rect 4486 1571 4546 1572
rect 2821 1545 2855 1571
rect 4512 1545 4546 1571
rect 2981 1504 3015 1520
rect 4355 1503 4389 1519
rect 2981 1409 3015 1470
rect 3227 1468 3243 1502
rect 3311 1468 3327 1502
rect 3499 1468 3515 1502
rect 3583 1468 3599 1502
rect 3771 1468 3787 1502
rect 3855 1468 3871 1502
rect 4043 1468 4059 1502
rect 4127 1468 4143 1502
rect 2981 1217 3015 1233
rect 3069 1409 3103 1425
rect 3069 1217 3103 1233
rect 3181 1409 3215 1425
rect 3181 1217 3215 1233
rect 3339 1409 3373 1425
rect 3339 1217 3373 1233
rect 3453 1409 3487 1425
rect 3453 1217 3487 1233
rect 3611 1409 3645 1425
rect 3611 1217 3645 1233
rect 3725 1409 3759 1425
rect 3725 1217 3759 1233
rect 3883 1409 3917 1425
rect 3883 1217 3917 1233
rect 3997 1409 4031 1425
rect 3997 1217 4031 1233
rect 4155 1409 4189 1425
rect 4155 1217 4189 1233
rect 4267 1409 4301 1425
rect 4267 1217 4301 1233
rect 4355 1409 4389 1469
rect 4355 1217 4389 1233
rect 3499 1140 3515 1174
rect 3583 1140 3599 1174
rect 3771 1140 3787 1174
rect 3855 1140 3871 1174
rect 3499 1032 3515 1066
rect 3583 1032 3599 1066
rect 3771 1032 3787 1066
rect 3855 1032 3871 1066
rect 2981 973 3015 989
rect 2981 726 3015 797
rect 3069 973 3103 989
rect 3069 781 3103 797
rect 3181 973 3215 989
rect 3181 781 3215 797
rect 3339 973 3373 989
rect 3339 781 3373 797
rect 3453 973 3487 989
rect 3453 781 3487 797
rect 3611 973 3645 989
rect 3611 781 3645 797
rect 3725 973 3759 989
rect 3725 781 3759 797
rect 3883 973 3917 989
rect 3883 781 3917 797
rect 3997 973 4031 989
rect 3997 781 4031 797
rect 4155 973 4189 989
rect 4155 781 4189 797
rect 4267 973 4301 989
rect 4267 781 4301 797
rect 4355 973 4389 989
rect 3227 704 3243 738
rect 3311 704 3327 738
rect 3499 704 3515 738
rect 3583 704 3599 738
rect 3771 704 3787 738
rect 3855 704 3871 738
rect 4043 704 4059 738
rect 4127 704 4143 738
rect 4355 734 4389 797
rect 2981 676 3015 692
rect 4355 684 4389 700
rect 2821 605 2855 631
rect 4512 606 4546 631
rect 2855 571 2881 605
rect 4486 571 4512 605
<< viali >>
rect 2803 1571 2855 1623
rect 4512 1572 4564 1624
rect 2981 1470 3015 1504
rect 3243 1468 3311 1502
rect 3515 1468 3583 1502
rect 3787 1468 3855 1502
rect 4059 1468 4127 1502
rect 4355 1469 4389 1503
rect 2981 1233 3015 1409
rect 3069 1233 3103 1409
rect 3181 1233 3215 1409
rect 3339 1233 3373 1409
rect 3453 1233 3487 1409
rect 3611 1233 3645 1409
rect 3725 1233 3759 1409
rect 3883 1233 3917 1409
rect 3997 1233 4031 1409
rect 4155 1233 4189 1409
rect 4267 1233 4301 1409
rect 4355 1233 4389 1409
rect 3515 1140 3583 1174
rect 3787 1140 3855 1174
rect 3515 1139 3583 1140
rect 3515 1032 3583 1066
rect 3787 1032 3855 1066
rect 2981 797 3015 973
rect 3069 797 3103 973
rect 3181 797 3215 973
rect 3339 797 3373 973
rect 3453 797 3487 973
rect 3611 797 3645 973
rect 3725 797 3759 973
rect 3883 797 3917 973
rect 3997 797 4031 973
rect 4155 797 4189 973
rect 4267 797 4301 973
rect 4355 797 4389 973
rect 2981 692 3015 726
rect 3243 704 3311 738
rect 3515 704 3583 738
rect 3787 704 3855 738
rect 4059 704 4127 738
rect 4355 700 4389 734
rect 2803 553 2855 605
rect 4512 554 4564 606
<< metal1 >>
rect 2791 1623 2867 1629
rect 2791 1571 2803 1623
rect 2855 1571 2867 1623
rect 4500 1624 4576 1630
rect 4500 1572 4512 1624
rect 4564 1572 4576 1624
rect 2791 1565 2867 1571
rect 2899 1567 3079 1571
rect 2899 1534 3102 1567
rect 2899 1223 2932 1534
rect 2975 1504 3021 1534
rect 2975 1470 2981 1504
rect 3015 1470 3021 1504
rect 2975 1409 3021 1470
rect 3069 1423 3102 1534
rect 3352 1538 4018 1567
rect 3231 1502 3323 1508
rect 3231 1468 3243 1502
rect 3311 1468 3323 1502
rect 3231 1462 3323 1468
rect 3069 1421 3205 1423
rect 3352 1421 3386 1538
rect 3503 1502 3595 1508
rect 3503 1468 3515 1502
rect 3583 1468 3595 1502
rect 3503 1462 3595 1468
rect 3665 1425 3705 1538
rect 3775 1502 3867 1508
rect 3775 1468 3787 1502
rect 3855 1468 3867 1502
rect 3775 1462 3867 1468
rect 2975 1233 2981 1409
rect 3015 1233 3021 1409
rect 2858 1159 2868 1223
rect 2932 1180 2942 1223
rect 2975 1221 3021 1233
rect 3063 1409 3221 1421
rect 3063 1233 3069 1409
rect 3103 1233 3181 1409
rect 3215 1233 3221 1409
rect 3063 1223 3221 1233
rect 3063 1221 3109 1223
rect 3175 1221 3221 1223
rect 3333 1409 3386 1421
rect 3333 1233 3339 1409
rect 3373 1233 3386 1409
rect 3447 1409 3493 1421
rect 3447 1349 3453 1409
rect 3333 1221 3386 1233
rect 3346 1217 3386 1221
rect 3417 1233 3453 1349
rect 3487 1349 3493 1409
rect 3604 1409 3765 1425
rect 3983 1422 4018 1538
rect 4267 1542 4470 1570
rect 4500 1566 4576 1572
rect 4047 1502 4139 1508
rect 4047 1468 4059 1502
rect 4127 1468 4139 1502
rect 4047 1462 4139 1468
rect 4267 1423 4300 1542
rect 3983 1421 4023 1422
rect 4170 1421 4300 1423
rect 4349 1512 4394 1542
rect 4349 1503 4395 1512
rect 4349 1469 4355 1503
rect 4389 1469 4395 1503
rect 4349 1454 4395 1469
rect 4349 1421 4394 1454
rect 3604 1397 3611 1409
rect 3487 1285 3497 1349
rect 3487 1233 3493 1285
rect 3417 1221 3493 1233
rect 3605 1233 3611 1397
rect 3645 1233 3725 1409
rect 3759 1233 3765 1409
rect 3877 1409 3923 1421
rect 3877 1359 3883 1409
rect 3870 1295 3883 1359
rect 3417 1180 3453 1221
rect 3605 1216 3765 1233
rect 3877 1233 3883 1295
rect 3917 1359 3923 1409
rect 3983 1409 4037 1421
rect 3917 1233 3955 1359
rect 3877 1221 3955 1233
rect 3514 1180 3524 1185
rect 2932 1159 3453 1180
rect 3503 1175 3524 1180
rect 2898 1144 3453 1159
rect 3498 1174 3524 1175
rect 3576 1180 3586 1185
rect 3576 1174 3595 1180
rect 3498 1140 3515 1174
rect 3503 1139 3515 1140
rect 3583 1139 3595 1174
rect 3503 1133 3524 1139
rect 3576 1133 3595 1139
rect 3513 1072 3523 1075
rect 3503 1067 3523 1072
rect 3499 1066 3523 1067
rect 3575 1072 3585 1075
rect 3575 1067 3595 1072
rect 3575 1066 3600 1067
rect 2901 1048 3453 1065
rect 2858 984 2868 1048
rect 2932 1025 3453 1048
rect 3499 1032 3515 1066
rect 3583 1032 3600 1066
rect 3503 1026 3523 1032
rect 2932 984 2942 1025
rect 3083 985 3202 986
rect 3413 985 3453 1025
rect 3513 1023 3523 1026
rect 3575 1026 3595 1032
rect 3575 1023 3585 1026
rect 3670 989 3702 1216
rect 3786 1180 3796 1183
rect 3775 1174 3796 1180
rect 3848 1180 3858 1183
rect 3917 1182 3955 1221
rect 3983 1233 3997 1409
rect 4031 1233 4037 1409
rect 3983 1221 4037 1233
rect 4149 1409 4307 1421
rect 4149 1233 4155 1409
rect 4189 1233 4267 1409
rect 4301 1233 4307 1409
rect 4149 1223 4307 1233
rect 4149 1221 4195 1223
rect 4261 1221 4307 1223
rect 4349 1409 4395 1421
rect 4349 1233 4355 1409
rect 4389 1233 4395 1409
rect 4349 1221 4395 1233
rect 4437 1222 4470 1542
rect 3983 1217 4023 1221
rect 4427 1182 4437 1222
rect 3848 1174 3867 1180
rect 3771 1140 3787 1174
rect 3855 1140 3872 1174
rect 3917 1158 4437 1182
rect 4501 1158 4511 1222
rect 3917 1144 4468 1158
rect 3771 1139 3796 1140
rect 3775 1134 3796 1139
rect 3786 1131 3796 1134
rect 3848 1139 3872 1140
rect 3848 1134 3867 1139
rect 3848 1131 3858 1134
rect 3784 1072 3794 1075
rect 3775 1067 3794 1072
rect 3771 1066 3794 1067
rect 3846 1072 3856 1075
rect 3846 1067 3867 1072
rect 3846 1066 3871 1067
rect 3771 1032 3787 1066
rect 3855 1032 3871 1066
rect 3775 1026 3794 1032
rect 3784 1023 3794 1026
rect 3846 1031 3871 1032
rect 3917 1048 4470 1068
rect 3846 1026 3867 1031
rect 3917 1027 4437 1048
rect 3846 1023 3856 1026
rect 3606 985 3763 989
rect 3917 985 3958 1027
rect 2900 643 2932 984
rect 2975 973 3021 985
rect 2975 797 2981 973
rect 3015 797 3021 973
rect 2975 785 3021 797
rect 3063 973 3221 985
rect 3063 797 3069 973
rect 3103 797 3181 973
rect 3215 797 3221 973
rect 3063 786 3221 797
rect 3063 785 3109 786
rect 3175 785 3221 786
rect 3333 982 3379 985
rect 3333 973 3382 982
rect 3333 797 3339 973
rect 3373 797 3382 973
rect 3413 973 3493 985
rect 3413 852 3453 973
rect 3333 785 3382 797
rect 3447 797 3453 852
rect 3487 916 3493 973
rect 3605 973 3765 985
rect 3487 852 3498 916
rect 3487 797 3493 852
rect 3447 785 3493 797
rect 3605 797 3611 973
rect 3645 797 3725 973
rect 3759 797 3765 973
rect 3877 973 3958 985
rect 3877 923 3883 973
rect 3873 843 3883 923
rect 3605 785 3765 797
rect 3877 797 3883 843
rect 3917 843 3958 973
rect 3988 973 4037 985
rect 3917 797 3923 843
rect 3877 785 3923 797
rect 3988 797 3997 973
rect 4031 797 4037 973
rect 3988 785 4037 797
rect 4149 973 4307 985
rect 4149 797 4155 973
rect 4189 797 4267 973
rect 4301 797 4307 973
rect 4149 785 4307 797
rect 4349 973 4395 985
rect 4427 984 4437 1027
rect 4501 984 4511 1048
rect 4349 797 4355 973
rect 4389 797 4395 973
rect 4349 785 4395 797
rect 2976 741 3021 785
rect 2975 726 3021 741
rect 2975 692 2981 726
rect 3015 692 3021 726
rect 2975 683 3021 692
rect 2976 643 3021 683
rect 3069 643 3102 785
rect 3335 781 3382 785
rect 3231 738 3323 744
rect 3231 704 3243 738
rect 3311 704 3323 738
rect 3231 698 3323 704
rect 2791 605 2867 611
rect 2900 610 3103 643
rect 3353 639 3382 781
rect 3503 738 3595 744
rect 3503 704 3515 738
rect 3583 704 3595 738
rect 3503 698 3595 704
rect 3665 639 3704 785
rect 3988 784 4035 785
rect 3775 738 3867 744
rect 3775 704 3787 738
rect 3855 704 3867 738
rect 3775 698 3867 704
rect 3989 639 4018 784
rect 4047 738 4139 744
rect 4047 704 4059 738
rect 4127 704 4139 738
rect 4047 698 4139 704
rect 3353 610 4018 639
rect 4267 643 4300 785
rect 4349 749 4394 785
rect 4349 734 4395 749
rect 4349 700 4355 734
rect 4389 700 4395 734
rect 4349 691 4395 700
rect 4349 643 4394 691
rect 4437 643 4470 984
rect 4267 610 4470 643
rect 2791 553 2803 605
rect 2855 553 2867 605
rect 2791 547 2867 553
rect 4500 606 4576 612
rect 4500 554 4512 606
rect 4564 554 4576 606
rect 4500 548 4576 554
<< via1 >>
rect 2868 1159 2932 1223
rect 3524 1174 3576 1185
rect 3524 1139 3576 1174
rect 3524 1133 3576 1139
rect 3523 1066 3575 1075
rect 2868 984 2932 1048
rect 3523 1032 3575 1066
rect 3523 1023 3575 1032
rect 3796 1174 3848 1183
rect 3796 1140 3848 1174
rect 4437 1158 4501 1222
rect 3796 1131 3848 1140
rect 3794 1066 3846 1075
rect 3794 1032 3846 1066
rect 3794 1023 3846 1032
rect 4437 984 4501 1048
<< metal2 >>
rect 2868 1223 2932 1233
rect 4416 1225 4521 1243
rect 2868 1149 2932 1159
rect 3522 1188 3578 1198
rect 3796 1184 3848 1193
rect 3522 1120 3578 1130
rect 3669 1183 3852 1184
rect 3669 1131 3796 1183
rect 3848 1131 3852 1183
rect 4416 1155 4433 1225
rect 4503 1155 4521 1225
rect 4416 1144 4521 1155
rect 3669 1130 3852 1131
rect 3523 1075 3575 1085
rect 3669 1075 3702 1130
rect 3796 1121 3848 1130
rect 2846 1050 2951 1064
rect 2846 980 2864 1050
rect 2929 1048 2951 1050
rect 2932 1047 2951 1048
rect 2934 980 2951 1047
rect 3522 1023 3523 1075
rect 3575 1023 3702 1075
rect 3522 1021 3702 1023
rect 3792 1078 3848 1088
rect 4437 1053 4501 1058
rect 3523 1013 3575 1021
rect 3792 1010 3848 1020
rect 4420 1048 4510 1053
rect 2846 965 2951 980
rect 4420 984 4437 1048
rect 4501 984 4510 1048
rect 4420 974 4510 984
<< via2 >>
rect 2868 1159 2932 1223
rect 3522 1185 3578 1188
rect 3522 1133 3524 1185
rect 3524 1133 3576 1185
rect 3576 1133 3578 1185
rect 3522 1130 3578 1133
rect 4433 1222 4503 1225
rect 4433 1158 4437 1222
rect 4437 1158 4501 1222
rect 4501 1158 4503 1222
rect 4433 1155 4503 1158
rect 2864 1048 2929 1050
rect 2864 984 2868 1048
rect 2868 1047 2929 1048
rect 2868 984 2932 1047
rect 2932 984 2934 1047
rect 2864 980 2934 984
rect 3792 1075 3848 1078
rect 3792 1023 3794 1075
rect 3794 1023 3846 1075
rect 3846 1023 3848 1075
rect 3792 1020 3848 1023
rect 4437 984 4501 1048
<< metal3 >>
rect 3111 1510 3988 1570
rect 2840 1227 2956 1243
rect 2840 1154 2862 1227
rect 2938 1154 2956 1227
rect 2840 1138 2956 1154
rect 3111 1072 3171 1510
rect 3928 1223 3988 1510
rect 4416 1225 4521 1243
rect 4416 1223 4433 1225
rect 3512 1188 3724 1193
rect 3512 1130 3522 1188
rect 3578 1130 3724 1188
rect 3928 1157 4433 1223
rect 3512 1124 3724 1130
rect 3645 1084 3724 1124
rect 3645 1078 3860 1084
rect 2895 1064 3443 1072
rect 2846 1050 3443 1064
rect 2846 980 2864 1050
rect 2929 1047 3443 1050
rect 2934 1012 3443 1047
rect 3645 1020 3792 1078
rect 3848 1020 3860 1078
rect 3645 1015 3860 1020
rect 3645 1014 3724 1015
rect 2934 980 2951 1012
rect 2846 965 2951 980
rect 3383 668 3443 1012
rect 4198 668 4258 1157
rect 4416 1155 4433 1157
rect 4503 1155 4521 1225
rect 4416 1144 4521 1155
rect 4414 1049 4519 1060
rect 4414 978 4432 1049
rect 4505 978 4519 1049
rect 4414 964 4519 978
rect 3383 608 4258 668
<< via3 >>
rect 2862 1223 2938 1227
rect 2862 1159 2868 1223
rect 2868 1159 2932 1223
rect 2932 1159 2938 1223
rect 2862 1154 2938 1159
rect 4432 1048 4505 1049
rect 4432 984 4437 1048
rect 4437 984 4501 1048
rect 4501 984 4505 1048
rect 4432 978 4505 984
<< metal4 >>
rect 3382 1508 4261 1568
rect 2840 1230 2956 1243
rect 3382 1230 3442 1508
rect 2840 1227 3442 1230
rect 2840 1154 2862 1227
rect 2938 1154 3442 1227
rect 2840 1151 3442 1154
rect 2840 1138 2956 1151
rect 3111 669 3171 1151
rect 4201 1060 4261 1508
rect 3927 1059 4519 1060
rect 3923 1049 4519 1059
rect 3923 980 4432 1049
rect 3923 669 3985 980
rect 4260 979 4432 980
rect 4414 978 4432 979
rect 4505 978 4519 1049
rect 4414 964 4519 978
rect 3111 609 3985 669
<< labels >>
flabel metal1 4572 1581 4572 1581 0 FreeSans 800 0 0 0 vdd
port 0 nsew
flabel metal2 3760 1146 3760 1146 0 FreeSans 800 0 0 0 vip
port 1 nsew
flabel metal3 3614 1152 3614 1152 0 FreeSans 800 0 0 0 vin
port 2 nsew
flabel metal1 3683 1453 3683 1453 0 FreeSans 800 0 0 0 d5
port 3 nsew
flabel metal4 3144 722 3144 722 0 FreeSans 800 0 0 0 d6
port 4 nsew
flabel metal3 4397 1195 4397 1195 0 FreeSans 800 0 0 0 out
port 5 nsew
<< end >>
