magic
tech sky130A
magscale 1 2
timestamp 1729222144
<< nmos >>
rect -80 527 80 727
rect -80 109 80 309
rect -80 -309 80 -109
rect -80 -727 80 -527
<< ndiff >>
rect -138 715 -80 727
rect -138 539 -126 715
rect -92 539 -80 715
rect -138 527 -80 539
rect 80 715 138 727
rect 80 539 92 715
rect 126 539 138 715
rect 80 527 138 539
rect -138 297 -80 309
rect -138 121 -126 297
rect -92 121 -80 297
rect -138 109 -80 121
rect 80 297 138 309
rect 80 121 92 297
rect 126 121 138 297
rect 80 109 138 121
rect -138 -121 -80 -109
rect -138 -297 -126 -121
rect -92 -297 -80 -121
rect -138 -309 -80 -297
rect 80 -121 138 -109
rect 80 -297 92 -121
rect 126 -297 138 -121
rect 80 -309 138 -297
rect -138 -539 -80 -527
rect -138 -715 -126 -539
rect -92 -715 -80 -539
rect -138 -727 -80 -715
rect 80 -539 138 -527
rect 80 -715 92 -539
rect 126 -715 138 -539
rect 80 -727 138 -715
<< ndiffc >>
rect -126 539 -92 715
rect 92 539 126 715
rect -126 121 -92 297
rect 92 121 126 297
rect -126 -297 -92 -121
rect 92 -297 126 -121
rect -126 -715 -92 -539
rect 92 -715 126 -539
<< poly >>
rect -80 799 80 815
rect -80 765 -64 799
rect 64 765 80 799
rect -80 727 80 765
rect -80 489 80 527
rect -80 455 -64 489
rect 64 455 80 489
rect -80 439 80 455
rect -80 381 80 397
rect -80 347 -64 381
rect 64 347 80 381
rect -80 309 80 347
rect -80 71 80 109
rect -80 37 -64 71
rect 64 37 80 71
rect -80 21 80 37
rect -80 -37 80 -21
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -80 -109 80 -71
rect -80 -347 80 -309
rect -80 -381 -64 -347
rect 64 -381 80 -347
rect -80 -397 80 -381
rect -80 -455 80 -439
rect -80 -489 -64 -455
rect 64 -489 80 -455
rect -80 -527 80 -489
rect -80 -765 80 -727
rect -80 -799 -64 -765
rect 64 -799 80 -765
rect -80 -815 80 -799
<< polycont >>
rect -64 765 64 799
rect -64 455 64 489
rect -64 347 64 381
rect -64 37 64 71
rect -64 -71 64 -37
rect -64 -381 64 -347
rect -64 -489 64 -455
rect -64 -799 64 -765
<< locali >>
rect -80 765 -64 799
rect 64 765 80 799
rect -126 715 -92 731
rect -126 523 -92 539
rect 92 715 126 731
rect 92 523 126 539
rect -80 455 -64 489
rect 64 455 80 489
rect -80 347 -64 381
rect 64 347 80 381
rect -126 297 -92 313
rect -126 105 -92 121
rect 92 297 126 313
rect 92 105 126 121
rect -80 37 -64 71
rect 64 37 80 71
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -126 -121 -92 -105
rect -126 -313 -92 -297
rect 92 -121 126 -105
rect 92 -313 126 -297
rect -80 -381 -64 -347
rect 64 -381 80 -347
rect -80 -489 -64 -455
rect 64 -489 80 -455
rect -126 -539 -92 -523
rect -126 -731 -92 -715
rect 92 -539 126 -523
rect 92 -731 126 -715
rect -80 -799 -64 -765
rect 64 -799 80 -765
<< viali >>
rect -64 765 64 799
rect -126 539 -92 715
rect 92 539 126 715
rect -64 455 64 489
rect -64 347 64 381
rect -126 121 -92 297
rect 92 121 126 297
rect -64 37 64 71
rect -64 -71 64 -37
rect -126 -297 -92 -121
rect 92 -297 126 -121
rect -64 -381 64 -347
rect -64 -489 64 -455
rect -126 -715 -92 -539
rect 92 -715 126 -539
rect -64 -799 64 -765
<< metal1 >>
rect -76 799 76 805
rect -76 765 -64 799
rect 64 765 76 799
rect -76 759 76 765
rect -132 715 -86 727
rect -132 539 -126 715
rect -92 539 -86 715
rect -132 527 -86 539
rect 86 715 132 727
rect 86 539 92 715
rect 126 539 132 715
rect 86 527 132 539
rect -76 489 76 495
rect -76 455 -64 489
rect 64 455 76 489
rect -76 449 76 455
rect -76 381 76 387
rect -76 347 -64 381
rect 64 347 76 381
rect -76 341 76 347
rect -132 297 -86 309
rect -132 121 -126 297
rect -92 121 -86 297
rect -132 109 -86 121
rect 86 297 132 309
rect 86 121 92 297
rect 126 121 132 297
rect 86 109 132 121
rect -76 71 76 77
rect -76 37 -64 71
rect 64 37 76 71
rect -76 31 76 37
rect -76 -37 76 -31
rect -76 -71 -64 -37
rect 64 -71 76 -37
rect -76 -77 76 -71
rect -132 -121 -86 -109
rect -132 -297 -126 -121
rect -92 -297 -86 -121
rect -132 -309 -86 -297
rect 86 -121 132 -109
rect 86 -297 92 -121
rect 126 -297 132 -121
rect 86 -309 132 -297
rect -76 -347 76 -341
rect -76 -381 -64 -347
rect 64 -381 76 -347
rect -76 -387 76 -381
rect -76 -455 76 -449
rect -76 -489 -64 -455
rect 64 -489 76 -455
rect -76 -495 76 -489
rect -132 -539 -86 -527
rect -132 -715 -126 -539
rect -92 -715 -86 -539
rect -132 -727 -86 -715
rect 86 -539 132 -527
rect 86 -715 92 -539
rect 126 -715 132 -539
rect 86 -727 132 -715
rect -76 -765 76 -759
rect -76 -799 -64 -765
rect 64 -799 76 -765
rect -76 -805 76 -799
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 4 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
