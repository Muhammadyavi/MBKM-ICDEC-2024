magic
tech sky130A
magscale 1 2
timestamp 1729216856
<< psubdiff >>
rect 974 572 1034 606
rect 2176 572 2236 606
rect 974 546 1008 572
rect 2202 546 2236 572
rect 974 -590 1008 -564
rect 2202 -590 2236 -564
rect 974 -624 1034 -590
rect 2176 -624 2236 -590
<< psubdiffcont >>
rect 1034 572 2176 606
rect 974 -564 1008 546
rect 2202 -564 2236 546
rect 1034 -624 2176 -590
<< poly >>
rect 1058 522 1207 538
rect 1058 488 1074 522
rect 1108 488 1162 522
rect 1196 488 1207 522
rect 1058 472 1207 488
rect 1520 478 1690 534
rect 2003 522 2152 538
rect 2003 488 2014 522
rect 2048 488 2102 522
rect 2136 488 2152 522
rect 2003 472 2152 488
rect 1120 446 1150 472
rect 2060 446 2090 472
rect 1520 -32 1690 14
rect 1120 -490 1150 -464
rect 2060 -486 2090 -460
rect 1058 -506 1207 -490
rect 1058 -540 1074 -506
rect 1108 -540 1162 -506
rect 1196 -540 1207 -506
rect 1058 -556 1207 -540
rect 1520 -552 1690 -497
rect 2003 -502 2152 -486
rect 2003 -536 2014 -502
rect 2048 -536 2102 -502
rect 2136 -536 2152 -502
rect 2003 -552 2152 -536
<< polycont >>
rect 1074 488 1108 522
rect 1162 488 1196 522
rect 2014 488 2048 522
rect 2102 488 2136 522
rect 1074 -540 1108 -506
rect 1162 -540 1196 -506
rect 2014 -536 2048 -502
rect 2102 -536 2136 -502
<< locali >>
rect 974 572 1034 606
rect 2176 572 2236 606
rect 974 546 1008 572
rect 2202 546 2236 572
rect 1074 522 1108 538
rect 1074 446 1108 488
rect 1162 522 1196 538
rect 1162 446 1196 488
rect 2014 522 2048 538
rect 2014 446 2048 488
rect 2102 522 2136 538
rect 2102 446 2136 488
rect 1074 -506 1108 -464
rect 1074 -556 1108 -540
rect 1162 -506 1196 -464
rect 1162 -556 1196 -540
rect 2014 -502 2048 -460
rect 2014 -552 2048 -536
rect 2102 -502 2136 -460
rect 2102 -552 2136 -536
rect 974 -590 1008 -564
rect 2202 -590 2236 -564
rect 974 -624 1034 -590
rect 2176 -624 2236 -590
<< viali >>
rect 1520 606 1578 616
rect 1520 572 1578 606
rect 1520 560 1578 572
rect 1074 488 1108 522
rect 1162 488 1196 522
rect 2014 488 2048 522
rect 2102 488 2136 522
rect 1074 -540 1108 -506
rect 1162 -540 1196 -506
rect 2014 -536 2048 -502
rect 2102 -536 2136 -502
rect 1633 -590 1689 -580
rect 1633 -624 1689 -590
rect 1633 -635 1689 -624
<< metal1 >>
rect 1508 616 1590 622
rect 1508 560 1520 616
rect 1578 560 1590 616
rect 1508 554 1590 560
rect 1068 522 1114 538
rect 1068 488 1074 522
rect 1108 488 1114 522
rect 1068 446 1114 488
rect 1156 522 1202 538
rect 1156 488 1162 522
rect 1196 488 1202 522
rect 1156 446 1202 488
rect 2008 522 2054 538
rect 2008 488 2014 522
rect 2048 488 2054 522
rect 2008 446 2054 488
rect 2096 522 2142 538
rect 2096 488 2102 522
rect 2136 488 2142 522
rect 2096 446 2142 488
rect 1179 64 1294 434
rect 1513 382 1523 434
rect 1575 382 1585 434
rect 1995 431 2005 434
rect 1911 382 2005 431
rect 2057 382 2067 434
rect 1179 58 1314 64
rect 1625 58 1635 110
rect 1687 58 1697 110
rect 1911 58 2026 382
rect 1268 14 1314 58
rect 1268 -32 1348 14
rect 1862 8 1942 14
rect 1858 -26 1942 8
rect 1862 -32 1942 -26
rect 1896 -64 1942 -32
rect 1178 -400 1294 -72
rect 1512 -128 1522 -76
rect 1574 -128 1584 -76
rect 1143 -452 1153 -400
rect 1205 -452 1294 -400
rect 1625 -452 1635 -400
rect 1687 -452 1697 -400
rect 1178 -454 1294 -452
rect 1919 -460 2031 -64
rect 1919 -462 2054 -460
rect 1068 -506 1114 -464
rect 1068 -540 1074 -506
rect 1108 -540 1114 -506
rect 1068 -556 1114 -540
rect 1156 -506 1202 -464
rect 1156 -540 1162 -506
rect 1196 -540 1202 -506
rect 1156 -556 1202 -540
rect 2008 -502 2054 -462
rect 2008 -536 2014 -502
rect 2048 -536 2054 -502
rect 2008 -552 2054 -536
rect 2096 -502 2142 -460
rect 2096 -536 2102 -502
rect 2136 -536 2142 -502
rect 2096 -552 2142 -536
rect 1621 -580 1701 -574
rect 1621 -636 1632 -580
rect 1690 -636 1701 -580
rect 1621 -641 1701 -636
<< via1 >>
rect 1520 560 1578 616
rect 1523 382 1575 434
rect 2005 382 2057 434
rect 1635 58 1687 110
rect 1522 -128 1574 -76
rect 1153 -452 1205 -400
rect 1635 -452 1687 -400
rect 1632 -635 1633 -580
rect 1633 -635 1689 -580
rect 1689 -635 1690 -580
rect 1632 -636 1690 -635
<< metal2 >>
rect 1520 616 1578 626
rect 1520 550 1578 560
rect 1521 436 1577 446
rect 1521 370 1577 380
rect 2001 438 2061 448
rect 2001 367 2061 377
rect 1635 110 1687 120
rect 1635 14 1687 58
rect 1522 -32 1687 14
rect 1522 -76 1574 -32
rect 1522 -138 1574 -128
rect 1148 -396 1210 -386
rect 1148 -466 1210 -456
rect 1633 -398 1689 -388
rect 1633 -464 1689 -454
rect 1149 -467 1209 -466
rect 1632 -580 1690 -570
rect 1632 -646 1690 -636
<< via2 >>
rect 1520 560 1578 616
rect 1521 434 1577 436
rect 1521 382 1523 434
rect 1523 382 1575 434
rect 1575 382 1577 434
rect 1521 380 1577 382
rect 2001 434 2061 438
rect 2001 382 2005 434
rect 2005 382 2057 434
rect 2057 382 2061 434
rect 2001 377 2061 382
rect 1148 -400 1210 -396
rect 1148 -452 1153 -400
rect 1153 -452 1205 -400
rect 1205 -452 1210 -400
rect 1148 -456 1210 -452
rect 1633 -400 1689 -398
rect 1633 -452 1635 -400
rect 1635 -452 1687 -400
rect 1687 -452 1689 -400
rect 1633 -454 1689 -452
rect 1632 -636 1690 -580
<< metal3 >>
rect 1507 616 1588 621
rect 1507 560 1520 616
rect 1578 560 1588 616
rect 1507 555 1588 560
rect 1507 447 1587 555
rect 1506 444 1589 447
rect 1506 436 1590 444
rect 1506 380 1521 436
rect 1577 380 1590 436
rect 1506 371 1590 380
rect 1964 441 2095 462
rect 1964 371 1995 441
rect 2066 371 2095 441
rect 1506 29 1589 371
rect 1964 347 2095 371
rect 1506 -47 1702 29
rect 1112 -392 1243 -373
rect 1112 -458 1145 -392
rect 1213 -458 1243 -392
rect 1112 -488 1243 -458
rect 1619 -398 1702 -47
rect 1619 -454 1633 -398
rect 1689 -454 1702 -398
rect 1619 -462 1702 -454
rect 1621 -580 1702 -462
rect 1621 -636 1632 -580
rect 1690 -636 1702 -580
rect 1621 -641 1702 -636
<< via3 >>
rect 1995 438 2066 441
rect 1995 377 2001 438
rect 2001 377 2061 438
rect 2061 377 2066 438
rect 1995 371 2066 377
rect 1145 -396 1213 -392
rect 1145 -456 1148 -396
rect 1148 -456 1210 -396
rect 1210 -456 1213 -396
rect 1145 -458 1213 -456
<< metal4 >>
rect 1977 441 2083 452
rect 1977 371 1995 441
rect 2066 371 2083 441
rect 1977 356 2083 371
rect 1995 25 2066 356
rect 1145 -42 2066 25
rect 1145 -379 1216 -42
rect 1127 -392 1233 -379
rect 1127 -458 1145 -392
rect 1213 -458 1233 -392
rect 1127 -475 1233 -458
use sky130_fd_pr__nfet_01v8_S44669  sky130_fd_pr__nfet_01v8_S44669_0
timestamp 1729216231
transform 1 0 1790 0 1 -264
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_S44669  sky130_fd_pr__nfet_01v8_S44669_2
timestamp 1729216231
transform 1 0 1420 0 1 246
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_S44669  sky130_fd_pr__nfet_01v8_S44669_3
timestamp 1729216231
transform 1 0 1790 0 1 246
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_S44669  sky130_fd_pr__nfet_01v8_S44669_4
timestamp 1729216231
transform 1 0 1420 0 1 -264
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_3
timestamp 1729182865
transform 1 0 1135 0 1 -264
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_5
timestamp 1729182865
transform 1 0 1135 0 1 246
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_6
timestamp 1729182865
transform 1 0 2075 0 1 246
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_7
timestamp 1729182865
transform 1 0 2075 0 1 -264
box -73 -226 73 226
<< labels >>
flabel space 1430 212 1430 212 0 FreeSans 320 0 0 0 m3
flabel space 1780 -392 1780 -392 0 FreeSans 320 0 0 0 m3
flabel space 1416 -390 1416 -390 0 FreeSans 320 0 0 0 m4
flabel space 1778 216 1778 216 0 FreeSans 320 0 0 0 m4
flabel space 1664 222 1664 222 0 FreeSans 320 0 0 0 rs
flabel space 1546 -390 1546 -390 0 FreeSans 320 0 0 0 rs
flabel metal2 1664 -390 1664 -390 0 FreeSans 320 0 0 0 s
flabel metal1 1286 -286 1286 -286 0 FreeSans 320 0 0 0 d4
flabel space 1916 -276 1916 -276 0 FreeSans 320 0 0 0 d3
flabel metal1 1290 221 1290 221 0 FreeSans 320 0 0 0 d3
flabel metal3 1548 226 1548 226 0 FreeSans 320 0 0 0 s
flabel metal1 1911 227 1911 227 0 FreeSans 320 0 0 0 d4
flabel metal4 2040 -24 2040 -24 0 FreeSans 640 0 0 0 d4
port 0 nsew
flabel metal2 1677 36 1677 36 0 FreeSans 640 0 0 0 rs
port 1 nsew
flabel metal1 1240 82 1240 82 0 FreeSans 640 0 0 0 d3
port 2 nsew
flabel metal3 1669 -480 1669 -480 0 FreeSans 640 0 0 0 gnd
port 3 nsew
<< end >>
