magic
tech sky130A
magscale 1 2
timestamp 1729337120
<< nwell >>
rect -1454 -575 -342 1682
rect -1454 -1792 1738 -575
<< viali >>
rect 1536 494 1676 634
rect 1537 299 1677 439
rect 1534 104 1674 244
rect 1538 -96 1678 44
rect 1538 -295 1678 -155
rect 1535 -495 1675 -355
<< metal1 >>
rect 1377 919 1387 1075
rect 1442 919 1452 1075
rect -271 816 6 850
rect -271 748 -237 816
rect -1397 594 -1387 677
rect -1309 650 -1299 677
rect -307 669 -297 748
rect -215 669 -205 748
rect -1309 610 -1161 650
rect -1309 594 -1299 610
rect -523 596 -513 663
rect -451 596 -441 663
rect -508 -1727 -472 -1293
rect -271 -1493 -237 669
rect 379 649 799 773
rect 1057 734 1674 770
rect 1562 640 1648 734
rect 1524 634 1688 640
rect -95 547 -85 614
rect 64 547 74 614
rect 1524 494 1536 634
rect 1676 494 1688 634
rect 1524 488 1688 494
rect 1525 439 1689 445
rect 1525 298 1536 439
rect 1677 298 1689 439
rect 1525 293 1689 298
rect 1522 248 1686 250
rect 1516 97 1526 248
rect 1684 97 1694 248
rect 1526 44 1690 50
rect 1526 -96 1538 44
rect 1678 -96 1690 44
rect 1526 -102 1690 -96
rect 1526 -150 1690 -149
rect 1516 -300 1526 -150
rect 1689 -300 1699 -150
rect 1526 -301 1690 -300
rect 1523 -355 1687 -349
rect -105 -482 -95 -415
rect -33 -482 -23 -415
rect 1523 -495 1535 -355
rect 1675 -495 1687 -355
rect 1523 -501 1687 -495
rect 1557 -647 1652 -501
rect -271 -1527 59 -1493
rect 711 -1727 747 -1323
rect 1137 -1474 1185 -1462
rect 1136 -1511 1185 -1474
rect 1137 -1695 1185 -1511
rect -508 -1763 747 -1727
rect 1110 -1767 1120 -1695
rect 1201 -1767 1211 -1695
<< via1 >>
rect 1387 919 1442 1075
rect -1387 594 -1309 677
rect -297 669 -215 748
rect -513 596 -451 663
rect -85 547 64 614
rect 1536 299 1537 439
rect 1537 299 1677 439
rect 1536 298 1677 299
rect 1526 244 1684 248
rect 1526 104 1534 244
rect 1534 104 1674 244
rect 1674 104 1684 244
rect 1526 97 1684 104
rect 1538 -96 1678 44
rect 1526 -155 1689 -150
rect 1526 -295 1538 -155
rect 1538 -295 1678 -155
rect 1678 -295 1689 -155
rect 1526 -300 1689 -295
rect -95 -482 -33 -415
rect 1120 -1767 1201 -1695
<< metal2 >>
rect 1380 1079 1447 1089
rect 1380 901 1447 911
rect -314 748 -201 762
rect -1386 687 -1308 688
rect -1397 678 -1299 687
rect -1397 677 -1386 678
rect -1397 594 -1387 677
rect -1397 593 -1386 594
rect -1308 593 -1299 678
rect -1397 585 -1299 593
rect -513 663 -451 673
rect -314 669 -297 748
rect -215 669 -201 748
rect -314 655 -201 669
rect 501 692 1141 726
rect -451 611 -343 648
rect -513 586 -451 596
rect -1387 584 -1308 585
rect -1386 583 -1308 584
rect -380 -430 -343 611
rect -85 614 64 624
rect -85 537 64 547
rect 501 131 535 692
rect 1107 187 1141 692
rect 1536 439 1677 449
rect 1536 288 1677 298
rect 1526 248 1684 258
rect 1107 153 1526 187
rect 1526 87 1684 97
rect 1538 44 1678 54
rect 1247 -60 1538 0
rect -95 -415 -33 -405
rect -380 -467 -95 -430
rect -95 -492 -33 -482
rect 1247 -1027 1307 -60
rect 1538 -106 1678 -96
rect 1526 -150 1689 -140
rect 1526 -310 1689 -300
rect 806 -1087 1307 -1027
rect 1103 -1695 1221 -1685
rect 1103 -1767 1120 -1695
rect 1201 -1767 1221 -1695
rect 1103 -1786 1221 -1767
<< via2 >>
rect 1380 1075 1447 1079
rect 1380 919 1387 1075
rect 1387 919 1442 1075
rect 1442 919 1447 1075
rect 1380 911 1447 919
rect -1386 677 -1308 678
rect -1387 594 -1309 677
rect -1309 594 -1308 677
rect -1386 593 -1308 594
rect -297 669 -215 748
rect -85 547 64 614
rect 1536 298 1677 439
rect 1526 -300 1689 -150
rect 1120 -1767 1201 -1695
<< metal3 >>
rect -1390 1527 -203 1599
rect -1390 687 -1318 1527
rect -275 1147 -203 1527
rect -275 1075 27 1147
rect -314 748 -201 762
rect -1397 683 -1299 687
rect -1397 678 -1298 683
rect -1397 677 -1386 678
rect -1397 594 -1387 677
rect -1397 593 -1386 594
rect -1308 593 -1298 678
rect -314 669 -297 748
rect -215 669 -201 748
rect -314 655 -201 669
rect -45 619 27 1075
rect 1370 1079 1457 1084
rect 1370 911 1380 1079
rect 1447 911 1457 1079
rect 1370 906 1457 911
rect -1397 588 -1298 593
rect -95 614 74 619
rect -1397 585 -1299 588
rect -95 547 -85 614
rect 64 547 74 614
rect -95 542 74 547
rect 1382 -545 1449 906
rect 1526 439 1687 444
rect 1526 298 1536 439
rect 1677 298 1687 439
rect 1526 293 1687 298
rect 1516 -150 1699 -145
rect 1516 -300 1526 -150
rect 1689 -300 1699 -150
rect 1516 -305 1699 -300
rect 1382 -612 1716 -545
rect 1649 -1170 1716 -612
rect 1485 -1237 1716 -1170
rect 1103 -1695 1221 -1685
rect 1103 -1767 1120 -1695
rect 1201 -1767 1221 -1695
rect 1103 -1786 1221 -1767
<< via3 >>
rect -297 669 -215 748
rect 1536 298 1677 439
rect 1526 -300 1689 -150
rect 1120 -1767 1201 -1695
<< metal4 >>
rect -314 748 -201 762
rect -314 669 -297 748
rect -215 742 -201 748
rect -215 674 1309 742
rect -215 669 -201 674
rect -314 655 -201 669
rect 1241 400 1309 674
rect 1535 439 1678 440
rect 1535 400 1536 439
rect 1241 332 1536 400
rect 1535 298 1536 332
rect 1677 298 1678 439
rect 1535 297 1678 298
rect 1525 -150 1690 -149
rect 1525 -199 1526 -150
rect 1130 -262 1526 -199
rect 1130 -487 1193 -262
rect 1525 -300 1526 -262
rect 1689 -300 1690 -150
rect 1525 -301 1690 -300
rect -241 -550 1193 -487
rect -241 -1700 -178 -550
rect 1103 -1695 1221 -1685
rect 1103 -1700 1120 -1695
rect -241 -1763 1120 -1700
rect 1103 -1767 1120 -1763
rect 1201 -1767 1221 -1695
rect 1103 -1786 1221 -1767
use nmosds2  nmosds2_0
timestamp 1729222144
transform 1 0 116 0 1 807
box -288 -72 1560 866
use nmosds  nmosds_0
timestamp 1729216856
transform 1 0 -1143 0 1 75
box 974 -646 2236 626
use pmoscs2  pmoscs2_0
timestamp 1729314602
transform 1 0 -2954 0 1 -2217
box 2785 535 4582 1641
use pmoscs  pmoscs_0
timestamp 1729157646
transform 1 0 -1158 0 1 -645
box -176 -811 822 2121
<< labels >>
flabel metal1 1682 -430 1682 -430 0 FreeSans 1120 0 0 0 vdd
port 0 nsew
flabel metal1 1687 -35 1687 -35 0 FreeSans 1120 0 0 0 vip
port 2 nsew
flabel via1 1677 165 1677 165 0 FreeSans 1120 0 0 0 rs
port 3 nsew
flabel metal1 1677 362 1677 362 0 FreeSans 1120 0 0 0 out
port 4 nsew
flabel metal1 1678 558 1678 558 0 FreeSans 1120 0 0 0 gnd
port 5 nsew
flabel via1 1687 -260 1687 -260 0 FreeSans 1120 0 0 0 vin
port 1 nsew
<< end >>
