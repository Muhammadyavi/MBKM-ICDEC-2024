magic
tech sky130A
magscale 1 2
timestamp 1729157646
<< nwell >>
rect -176 -811 822 2121
<< nsubdiff >>
rect -140 2051 -80 2085
rect 726 2051 786 2085
rect -140 2013 -106 2051
rect 752 2013 786 2051
rect -140 -741 -106 -715
rect 752 -741 786 -715
rect -140 -775 -80 -741
rect 726 -775 786 -741
<< nsubdiffcont >>
rect -80 2051 726 2085
rect -140 -715 -106 2013
rect 752 -715 786 2013
rect -80 -775 726 -741
<< poly >>
rect -56 2001 36 2017
rect -56 1967 -40 2001
rect -6 1967 36 2001
rect -56 1951 36 1967
rect 6 1920 36 1951
rect 610 2001 702 2017
rect 610 1967 652 2001
rect 686 1967 702 2001
rect 610 1951 702 1967
rect 610 1920 640 1951
rect 94 1307 294 1423
rect -56 1291 36 1307
rect -56 1257 -40 1291
rect -6 1257 36 1291
rect -56 1241 36 1257
rect 6 1210 36 1241
rect 610 1291 702 1307
rect 610 1257 652 1291
rect 686 1257 702 1291
rect 610 1241 702 1257
rect 610 1210 640 1241
rect 94 597 552 713
rect 6 69 36 100
rect -56 53 36 69
rect -56 19 -40 53
rect -6 19 36 53
rect -56 3 36 19
rect 610 69 640 100
rect 610 53 702 69
rect 610 19 652 53
rect 686 19 702 53
rect 610 3 702 19
rect 352 -113 552 3
rect 6 -641 36 -610
rect -56 -657 36 -641
rect -56 -691 -40 -657
rect -6 -691 36 -657
rect -56 -707 36 -691
rect 610 -641 640 -614
rect 610 -657 702 -641
rect 610 -691 652 -657
rect 686 -691 702 -657
rect 610 -707 702 -691
<< polycont >>
rect -40 1967 -6 2001
rect 652 1967 686 2001
rect -40 1257 -6 1291
rect 652 1257 686 1291
rect -40 19 -6 53
rect 652 19 686 53
rect -40 -691 -6 -657
rect 652 -691 686 -657
<< locali >>
rect -140 2051 -80 2085
rect 726 2051 786 2085
rect -140 2013 -106 2051
rect -40 2001 -6 2017
rect -40 1920 -6 1967
rect 652 2001 686 2017
rect 652 1920 686 1967
rect 752 2013 786 2051
rect -40 1291 -6 1307
rect -40 1210 -6 1257
rect 652 1291 686 1307
rect 652 1210 686 1257
rect -40 53 -6 100
rect -40 3 -6 19
rect 652 53 686 100
rect 652 3 686 19
rect -40 -657 -6 -610
rect -40 -707 -6 -691
rect 652 -657 686 -610
rect 652 -707 686 -691
rect -140 -741 -106 -715
rect 752 -741 786 -715
rect -140 -775 -80 -741
rect 726 -775 786 -741
<< viali >>
rect -40 1967 -6 2001
rect 652 1967 686 2001
rect 752 1967 786 2001
rect -40 1257 -6 1291
rect 652 1257 686 1291
rect -40 19 -6 53
rect 652 19 686 53
rect -140 -691 -106 -657
rect -40 -691 -6 -657
rect 652 -691 686 -657
<< metal1 >>
rect -46 2001 0 2013
rect -46 1967 -40 2001
rect -6 1967 0 2001
rect -46 1920 0 1967
rect 646 2007 692 2013
rect 646 2001 798 2007
rect 646 1967 652 2001
rect 686 1967 752 2001
rect 786 1967 798 2001
rect 646 1961 798 1967
rect 646 1921 692 1961
rect 558 1920 692 1921
rect -46 1908 87 1920
rect -59 1532 -49 1908
rect 3 1532 87 1908
rect -49 1520 87 1532
rect -49 1445 3 1520
rect 299 1478 346 1920
rect 558 1908 691 1920
rect 558 1532 643 1908
rect 695 1532 705 1908
rect 558 1521 695 1532
rect 560 1478 606 1521
rect -59 1393 -49 1445
rect 3 1393 13 1445
rect 299 1432 606 1478
rect 645 1465 695 1521
rect 644 1445 696 1465
rect -46 1291 0 1303
rect -46 1257 -40 1291
rect -6 1257 0 1291
rect -46 1210 0 1257
rect -46 1198 87 1210
rect -46 822 39 1198
rect 91 822 101 1198
rect -46 810 87 822
rect 39 547 194 581
rect 39 500 92 547
rect -46 488 92 500
rect -59 487 92 488
rect -59 112 39 487
rect -46 111 39 112
rect 92 111 102 487
rect -46 100 87 111
rect -46 53 0 100
rect -46 19 -40 53
rect -6 19 0 53
rect -46 7 0 19
rect -60 -123 -50 -71
rect 2 -123 12 -71
rect 299 -122 346 1432
rect 634 1393 644 1445
rect 696 1393 706 1445
rect 646 1291 692 1303
rect 646 1257 652 1291
rect 686 1257 692 1291
rect 646 1210 692 1257
rect 559 1198 692 1210
rect 545 822 555 1198
rect 608 822 705 1198
rect 555 810 692 822
rect 555 763 608 810
rect 453 729 608 763
rect 559 488 692 500
rect 545 112 555 488
rect 607 112 692 488
rect 559 100 692 112
rect 646 53 692 100
rect 646 19 652 53
rect 686 19 692 53
rect 646 7 692 19
rect -50 -210 2 -123
rect 41 -169 346 -122
rect 632 -123 642 -71
rect 694 -123 704 -71
rect 41 -210 88 -169
rect -50 -222 88 -210
rect -60 -598 -50 -222
rect 2 -598 88 -222
rect -45 -610 88 -598
rect 299 -610 346 -169
rect 642 -210 694 -123
rect 558 -222 694 -210
rect 558 -598 642 -222
rect 694 -598 704 -222
rect 558 -610 692 -598
rect -46 -651 0 -610
rect -152 -657 0 -651
rect -152 -691 -140 -657
rect -106 -691 -40 -657
rect -6 -691 0 -657
rect -152 -697 0 -691
rect -46 -703 0 -697
rect 646 -657 692 -610
rect 646 -691 652 -657
rect 686 -691 692 -657
rect 646 -703 692 -691
<< via1 >>
rect -49 1532 3 1908
rect 643 1532 695 1908
rect -49 1393 3 1445
rect 39 822 91 1198
rect 39 111 92 487
rect -50 -123 2 -71
rect 644 1393 696 1445
rect 555 822 608 1198
rect 555 112 607 488
rect 642 -123 694 -71
rect -50 -598 2 -222
rect 642 -598 694 -222
<< metal2 >>
rect -49 1908 3 1918
rect -50 1532 -49 1533
rect 643 1908 695 1918
rect -50 1457 3 1532
rect 642 1532 643 1551
rect 642 1465 695 1532
rect 642 1457 696 1465
rect -51 1447 5 1457
rect -51 1381 5 1391
rect 642 1447 698 1457
rect 642 1381 698 1391
rect 39 1198 91 1208
rect 39 681 91 822
rect 555 1198 608 1208
rect 555 812 608 822
rect 39 629 607 681
rect 39 487 92 497
rect 39 101 92 111
rect 555 488 607 629
rect 555 102 607 112
rect -52 -69 4 -59
rect -52 -222 4 -125
rect 640 -69 696 -59
rect 640 -135 696 -125
rect -52 -226 -50 -222
rect 2 -226 4 -222
rect 642 -143 695 -135
rect 642 -222 694 -143
rect -50 -608 2 -598
rect 642 -608 694 -598
<< via2 >>
rect -51 1445 5 1447
rect -51 1393 -49 1445
rect -49 1393 3 1445
rect 3 1393 5 1445
rect -51 1391 5 1393
rect 642 1445 698 1447
rect 642 1393 644 1445
rect 644 1393 696 1445
rect 696 1393 698 1445
rect 642 1391 698 1393
rect -52 -71 4 -69
rect -52 -123 -50 -71
rect -50 -123 2 -71
rect 2 -123 4 -71
rect -52 -125 4 -123
rect 640 -71 696 -69
rect 640 -123 642 -71
rect 642 -123 694 -71
rect 694 -123 696 -71
rect 640 -125 696 -123
<< metal3 >>
rect -79 1447 29 1465
rect -79 1391 -51 1447
rect 5 1391 29 1447
rect -79 1366 29 1391
rect 614 1447 722 1465
rect 614 1391 642 1447
rect 698 1391 722 1447
rect 614 1367 722 1391
rect -55 686 8 1366
rect 281 746 291 810
rect 355 809 365 810
rect 640 809 703 1367
rect 355 746 703 809
rect -55 623 700 686
rect -52 500 291 563
rect -52 -45 11 500
rect 281 499 291 500
rect 355 499 365 563
rect 637 -44 700 623
rect -76 -69 32 -45
rect -76 -125 -52 -69
rect 4 -125 32 -69
rect -76 -143 32 -125
rect 616 -69 724 -44
rect 616 -125 640 -69
rect 696 -125 724 -69
rect 616 -143 724 -125
<< via3 >>
rect 291 746 355 810
rect 291 499 355 563
<< metal4 >>
rect 285 810 360 814
rect 285 746 291 810
rect 355 746 360 810
rect 285 563 360 746
rect 285 499 291 563
rect 355 499 360 563
rect 285 492 360 499
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_0
timestamp 1729132709
transform 1 0 625 0 1 -410
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_1
timestamp 1729132709
transform 1 0 21 0 1 1010
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_2
timestamp 1729132709
transform 1 0 21 0 1 -410
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_3
timestamp 1729132709
transform 1 0 21 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_4
timestamp 1729132709
transform 1 0 625 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_5
timestamp 1729132709
transform 1 0 625 0 1 1010
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_6
timestamp 1729132709
transform 1 0 21 0 1 1720
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_7
timestamp 1729132709
transform 1 0 625 0 1 1720
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729141416
transform 1 0 323 0 1 1720
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729141416
transform 1 0 323 0 1 1010
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729141416
transform 1 0 323 0 1 300
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729141416
transform 1 0 323 0 1 -410
box -323 -300 323 300
<< labels >>
flabel metal3 669 647 669 647 0 FreeSans 480 0 0 0 d5
port 0 nsew
flabel metal2 64 730 64 730 0 FreeSans 480 0 0 0 d1
port 1 nsew
flabel metal1 575 733 575 733 0 FreeSans 480 0 0 0 d2
port 2 nsew
flabel metal1 585 1490 585 1490 0 FreeSans 480 0 0 0 vdd
port 3 nsew
<< end >>
