magic
tech sky130A
magscale 1 2
timestamp 1729225416
<< error_p >>
rect -381 18 381 236
<< nwell >>
rect -381 18 381 418
rect -381 -418 381 -18
<< pmos >>
rect -287 118 -187 318
rect -129 118 -29 318
rect 29 118 129 318
rect 187 118 287 318
rect -287 -318 -187 -118
rect -129 -318 -29 -118
rect 29 -318 129 -118
rect 187 -318 287 -118
<< pdiff >>
rect -345 306 -287 318
rect -345 130 -333 306
rect -299 130 -287 306
rect -345 118 -287 130
rect -187 306 -129 318
rect -187 130 -175 306
rect -141 130 -129 306
rect -187 118 -129 130
rect -29 306 29 318
rect -29 130 -17 306
rect 17 130 29 306
rect -29 118 29 130
rect 129 306 187 318
rect 129 130 141 306
rect 175 130 187 306
rect 129 118 187 130
rect 287 306 345 318
rect 287 130 299 306
rect 333 130 345 306
rect 287 118 345 130
rect -345 -130 -287 -118
rect -345 -306 -333 -130
rect -299 -306 -287 -130
rect -345 -318 -287 -306
rect -187 -130 -129 -118
rect -187 -306 -175 -130
rect -141 -306 -129 -130
rect -187 -318 -129 -306
rect -29 -130 29 -118
rect -29 -306 -17 -130
rect 17 -306 29 -130
rect -29 -318 29 -306
rect 129 -130 187 -118
rect 129 -306 141 -130
rect 175 -306 187 -130
rect 129 -318 187 -306
rect 287 -130 345 -118
rect 287 -306 299 -130
rect 333 -306 345 -130
rect 287 -318 345 -306
<< pdiffc >>
rect -333 130 -299 306
rect -175 130 -141 306
rect -17 130 17 306
rect 141 130 175 306
rect 299 130 333 306
rect -333 -306 -299 -130
rect -175 -306 -141 -130
rect -17 -306 17 -130
rect 141 -306 175 -130
rect 299 -306 333 -130
<< poly >>
rect -287 399 -187 415
rect -287 365 -271 399
rect -203 365 -187 399
rect -287 318 -187 365
rect -129 399 -29 415
rect -129 365 -113 399
rect -45 365 -29 399
rect -129 318 -29 365
rect 29 399 129 415
rect 29 365 45 399
rect 113 365 129 399
rect 29 318 129 365
rect 187 399 287 415
rect 187 365 203 399
rect 271 365 287 399
rect 187 318 287 365
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -118 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -118 287 -71
rect -287 -365 -187 -318
rect -287 -399 -271 -365
rect -203 -399 -187 -365
rect -287 -415 -187 -399
rect -129 -365 -29 -318
rect -129 -399 -113 -365
rect -45 -399 -29 -365
rect -129 -415 -29 -399
rect 29 -365 129 -318
rect 29 -399 45 -365
rect 113 -399 129 -365
rect 29 -415 129 -399
rect 187 -365 287 -318
rect 187 -399 203 -365
rect 271 -399 287 -365
rect 187 -415 287 -399
<< polycont >>
rect -271 365 -203 399
rect -113 365 -45 399
rect 45 365 113 399
rect 203 365 271 399
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect -271 -399 -203 -365
rect -113 -399 -45 -365
rect 45 -399 113 -365
rect 203 -399 271 -365
<< locali >>
rect -287 365 -271 399
rect -203 365 -187 399
rect -129 365 -113 399
rect -45 365 -29 399
rect 29 365 45 399
rect 113 365 129 399
rect 187 365 203 399
rect 271 365 287 399
rect -333 306 -299 322
rect -333 114 -299 130
rect -175 306 -141 322
rect -175 114 -141 130
rect -17 306 17 322
rect -17 114 17 130
rect 141 306 175 322
rect 141 114 175 130
rect 299 306 333 322
rect 299 114 333 130
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect -333 -130 -299 -114
rect -333 -322 -299 -306
rect -175 -130 -141 -114
rect -175 -322 -141 -306
rect -17 -130 17 -114
rect -17 -322 17 -306
rect 141 -130 175 -114
rect 141 -322 175 -306
rect 299 -130 333 -114
rect 299 -322 333 -306
rect -287 -399 -271 -365
rect -203 -399 -187 -365
rect -129 -399 -113 -365
rect -45 -399 -29 -365
rect 29 -399 45 -365
rect 113 -399 129 -365
rect 187 -399 203 -365
rect 271 -399 287 -365
<< viali >>
rect -271 365 -203 399
rect -113 365 -45 399
rect 45 365 113 399
rect 203 365 271 399
rect -333 130 -299 306
rect -175 130 -141 306
rect -17 130 17 306
rect 141 130 175 306
rect 299 130 333 306
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect -333 -306 -299 -130
rect -175 -306 -141 -130
rect -17 -306 17 -130
rect 141 -306 175 -130
rect 299 -306 333 -130
rect -271 -399 -203 -365
rect -113 -399 -45 -365
rect 45 -399 113 -365
rect 203 -399 271 -365
<< metal1 >>
rect -283 399 -191 405
rect -283 365 -271 399
rect -203 365 -191 399
rect -283 359 -191 365
rect -125 399 -33 405
rect -125 365 -113 399
rect -45 365 -33 399
rect -125 359 -33 365
rect 33 399 125 405
rect 33 365 45 399
rect 113 365 125 399
rect 33 359 125 365
rect 191 399 283 405
rect 191 365 203 399
rect 271 365 283 399
rect 191 359 283 365
rect -339 306 -293 318
rect -339 130 -333 306
rect -299 130 -293 306
rect -339 118 -293 130
rect -181 306 -135 318
rect -181 130 -175 306
rect -141 130 -135 306
rect -181 118 -135 130
rect -23 306 23 318
rect -23 130 -17 306
rect 17 130 23 306
rect -23 118 23 130
rect 135 306 181 318
rect 135 130 141 306
rect 175 130 181 306
rect 135 118 181 130
rect 293 306 339 318
rect 293 130 299 306
rect 333 130 339 306
rect 293 118 339 130
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect -339 -130 -293 -118
rect -339 -306 -333 -130
rect -299 -306 -293 -130
rect -339 -318 -293 -306
rect -181 -130 -135 -118
rect -181 -306 -175 -130
rect -141 -306 -135 -130
rect -181 -318 -135 -306
rect -23 -130 23 -118
rect -23 -306 -17 -130
rect 17 -306 23 -130
rect -23 -318 23 -306
rect 135 -130 181 -118
rect 135 -306 141 -130
rect 175 -306 181 -130
rect 135 -318 181 -306
rect 293 -130 339 -118
rect 293 -306 299 -130
rect 333 -306 339 -130
rect 293 -318 339 -306
rect -283 -365 -191 -359
rect -283 -399 -271 -365
rect -203 -399 -191 -365
rect -283 -405 -191 -399
rect -125 -365 -33 -359
rect -125 -399 -113 -365
rect -45 -399 -33 -365
rect -125 -405 -33 -399
rect 33 -365 125 -359
rect 33 -399 45 -365
rect 113 -399 125 -365
rect 33 -405 125 -399
rect 191 -365 283 -359
rect 191 -399 203 -365
rect 271 -399 283 -365
rect 191 -405 283 -399
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
